
package aes_pkg;

  import uvm_pkg::*;
  typedef uvm_config_db#(virtual aes_interface) aes_vif_config;

  `include "uvm_macros.svh" 
  `include "aes_packet.sv"

  `include "aes_monitor.sv"
  `include "aes_monitor2.sv"
  `include "aes_sequencer.sv"
  `include "aes_seqs.sv"
  `include "aes_driver.sv"
  `include "aes_agent.sv"
  `include "aes_agent2.sv"
  `include "aes_env.sv" 
 

endpackage
